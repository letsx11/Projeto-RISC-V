`timescale 1ns / 1ps

module flopr #(
    parameter WIDTH = 8
) (
    input  logic clk,
    input  logic reset,
    input  logic [WIDTH-1:0] d,
    input  logic stall,
    input  logic halt,                  
    output logic [WIDTH-1:0] q
);

    always_ff @(posedge clk) begin
        if (reset)
            q <= 0;

        else if (halt)
            q <= q;                     

        else if (!stall)
            q <= d;
    end

endmodule
